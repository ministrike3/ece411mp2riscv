module pick_the_word 
(
input logic x
);
endmodule